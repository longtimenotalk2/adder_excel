.inc '/ic/projects/BM1374/public/5_custom/release/stdcell/stdcell_BM/elvt/spf/Cbest45/INVD1BM156H3P48CPDELVT_1.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/stdcell/stdcell_BM/elvt/spf/Cbest45/ND2D1BM156H3P48CPDELVT_1.Cbest45.spf'
.inc '/ic/projects/BM1374/users/haiwei.li/V0/work/spf/out/ND2D1BM156H3P48CPDELVT_1_H2H_V03/ND2D1BM156H3P48CPDELVT_1_H2H_V03.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/stdcell/stdcell_BM/elvt/spf/Cbest45/NR2D1BM156H3P48CPDELVT_1.Cbest45.spf'
.inc '/ic/projects/BM1374/users/haiwei.li/V0/work/spf/out/NR2D1BM156H3P48CPDELVT_1_H2H_V02/NR2D1BM156H3P48CPDELVT_1_H2H_V02.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/stdcell/stdcell_BM/elvt/spf/Cbest45/OR2D1BM156H3P48CPDELVT_1.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/stdcell/stdcell_BM/elvt/spf/Cbest45/IND2D1BM156H3P48CPDELVT_1.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/custom/elvt/spf/Cbest45/XOR2D1BM156H3P48CPDELVT.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/custom/elvt/spf/Cbest45/XNR2D1BM156H3P48CPDELVT.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/custom/elvt/spf/Cbest45/XOR2D1_DUAL_OUT_BM156H3P48CPDELVT.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/custom/elvt/spf/Cbest45/XNR2D1_DUAL_OUT_BM156H3P48CPDELVT.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/custom/elvt/spf/Cbest45/AOI21D1BM156H3P48CPDELVT.Cbest45.spf'
.inc '/ic/projects/BM1374/users/haiwei.li/V0/work/spf/out/AOI21D1BM156H3P48CPDELVT_H2H_V03/AOI21D1BM156H3P48CPDELVT_H2H_V03.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/custom/elvt/spf/Cbest45/AOI21D2BM156H3P48CPDELVT.Cbest45.spf'
.inc '/ic/projects/BM1374/users/haiwei.li/V0/work/spf/out/AOI21D2BM156H3P48CPDELVT_H2H_V03/AOI21D2BM156H3P48CPDELVT_H2H_V03.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/custom/elvt/spf/Cbest45/OAI21D1BM156H3P48CPDELVT.Cbest45.spf'
.inc '/ic/projects/BM1374/users/haiwei.li/V0/work/spf/out/OAI21D1BM156H3P48CPDELVT_H2H_V02/OAI21D1BM156H3P48CPDELVT_H2H_V02.Cbest45.spf'
.inc '/ic/projects/BM1374/users/haiwei.li/V0/work/spf/out/OAI21D2BM156H3P48CPDELVT_H2H_V02/OAI21D2BM156H3P48CPDELVT_H2H_V02.Cbest45.spf'
.inc '/ic/projects/BM1374/users/haiwei.li/V0/work/spf/out/OAI21D2BM156H3P48CPDELVT_H2H_V02/OAI21D2BM156H3P48CPDELVT_H2H_V02.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/custom/elvt/spf/Cbest45/OA21D1BM156H3P48CPDELVT.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/custom/elvt/spf/Cbest45/IAOI21D1BM156H3P48CPDELVT.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/custom/elvt/spf/Cbest45/AOI22D1BM156H3P48CPDELVT.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/stdcell/stdcell_BM/elvt/spf/Cbest45/AOI22D2BM156H3P48CPDELVT_1.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/custom/elvt/spf/Cbest45/OAI22D1BM156H3P48CPDELVT.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/custom/elvt/spf/Cbest45/OAOI211D1BM156H3P48CPDELVT.Cbest45.spf'
.inc '/ic/projects/BM1374/public/5_custom/release/custom/elvt/spf/Cbest45/OAO211D1BM156H3P48CPDELVT.Cbest45.spf'

.inc 'cell/hack_OAI22D1BM156H3P48CPDELVT_P_ULVTLL_L2H_V02.Cbest45.spf'
.inc 'cell/hack_OAI22D2BM156H3P48CPDELVT_1_P_ULVTLL_L2H.Cbest45.spf'
.inc 'cell/hack_NR2D1BM156H3P48CPDELVT_1_P_ULVTLL_L2H_V02.Cbest45.spf'

.SUBCKT VDH_UFADDER_PN_B04_T01 A0 A1 A2 A3 A4 A5 A6 A7 A8 A9 A10 A11 A12 A13 A14 A15 A16 A17 A18 A19 A20 A21 A22 A23 A24 A25 A26 A27 A28 A29 A30 B0 B1 B2 B3 B4 B5 B6 B7 B8 B9 B10 B11 B12 B13 B14 B15 B16 B17 B18 B19 B20 B21 B22 B23 B24 B25 B26 B27 B28 B29 B30 S0 S1 S2 S3 S4 S5 S6 S7 S8 S9 S10 S11 S12 S13 S14 S15 S16 S17 S18 S19 S20 S21 S22 S23 S24 S25 S26 S27 S28 S29 S30 VBB VDD VDDH VPP VSS 
x_U1_nh1_0          a1      b1      a0      b0      VBB     VDD     VPP     VSS     nh1_0    AOI22D2BM156H3P48CPDELVT_1
x_U1_np2_1          a2      b2      a1      b1      VBB     VDD     VPP     VSS     np2_1    OAI22D1BM156H3P48CPDELVT
x_U1_nh3_2          a3      b3      a2      b2      VBB     VDD     VPP     VSS     nh3_2    AOI22D2BM156H3P48CPDELVT_1
x_U1_np4_3          a4      b4      a3      b3      VBB     VDD     VPP     VSS     np4_3    OAI22D1BM156H3P48CPDELVT
x_U1_nh5_4          a5      b5      a4      b4      VBB     VDD     VPP     VSS     nh5_4    AOI22D1BM156H3P48CPDELVT
x_U1_np6_5          a6      b6      a5      b5      VBB     VDD     VPP     VSS     np6_5    OAI22D1BM156H3P48CPDELVT
x_U1_nh7_6          a7      b7      a6      b6      VBB     VDD     VPP     VSS     nh7_6    AOI22D1BM156H3P48CPDELVT
x_U1_np8_7          a8      b8      a7      b7      VBB     VDD     VPP     VSS     np8_7    OAI22D1BM156H3P48CPDELVT
x_U1_nh9_8          a9      b9      a8      b8      VBB     VDD     VPP     VSS     nh9_8    AOI22D1BM156H3P48CPDELVT
x_U1_np10_9         a10     b10     a9      b9      VBB     VDD     VPP     VSS     np10_9    OAI22D1BM156H3P48CPDELVT
x_U1_nh11_10        a11     b11     a10     b10     VBB     VDD     VPP     VSS     nh11_10    AOI22D1BM156H3P48CPDELVT
x_U1_np12_11        a12     b12     a11     b11     VBB     VDD     VPP     VSS     np12_11    OAI22D1BM156H3P48CPDELVT
x_U1_nh13_12        a13     b13     a12     b12     VBB     VDD     VPP     VSS     nh13_12    AOI22D1BM156H3P48CPDELVT
x_U1_np14_13        a14     b14     a13     b13     VBB     VDD     VPP     VSS     np14_13    OAI22D1BM156H3P48CPDELVT
x_U1_nh15_14        a15     b15     a14     b14     VBB     VDD     VPP     VSS     nh15_14    AOI22D1BM156H3P48CPDELVT
x_U1_np16_15        a16     b16     a15     b15     VBB     VDD     VPP     VSS     np16_15    OAI22D1BM156H3P48CPDELVT
x_U1_nh17_16        a17     b17     a16     b16     VBB     VDD     VPP     VSS     nh17_16    AOI22D1BM156H3P48CPDELVT
x_U1_np18_17        a18     b18     a17     b17     VBB     VDD     VPP     VSS     np18_17    OAI22D1BM156H3P48CPDELVT
x_U1_nh19_18        a19     b19     a18     b18     VBB     VDD     VPP     VSS     nh19_18    AOI22D1BM156H3P48CPDELVT
x_U1_np20_19        a20     b20     a19     b19     VBB     VDD     VPP     VSS     np20_19    OAI22D1BM156H3P48CPDELVT
x_U1_nh21_20        a21     b21     a20     b20     VBB     VDD     VPP     VSS     nh21_20    AOI22D1BM156H3P48CPDELVT
x_U1_np22_21        a22     b22     a21     b21     VBB     VDD     VPP     VSS     np22_21    OAI22D1BM156H3P48CPDELVT
x_U1_nh23_22        a23     b23     a22     b22     VBB     VDD     VPP     VSS     nh23_22    AOI22D1BM156H3P48CPDELVT
x_U1_np24_23        a24     b24     a23     b23     VBB     VDD     VPP     VSS     np24_23    OAI22D1BM156H3P48CPDELVT
x_U1_nh25_24        a25     b25     a24     b24     VBB     VDD     VPP     VSS     nh25_24    AOI22D1BM156H3P48CPDELVT
x_U1_np26_25        a26     b26     a25     b25     VBB     VDD     VPP     VSS     np26_25    OAI22D1BM156H3P48CPDELVT
x_U1_nh27_26        a27     b27     a26     b26     VBB     VDD     VPP     VSS     nh27_26    AOI22D1BM156H3P48CPDELVT
x_U1_np27_q27       a27     b27     np27    VBB     VDD     VPP     VSS     q27     XOR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_np28_q28       a28     b28     np28    VBB     VDD     VPP     VSS     q28     XOR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_ng29_nq29      a29     b29     ng29    VBB     VDD     VPP     VSS     nq29    XNR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U2_h3_0           np2_1    nh1_0    nh3_2    nh3_2    VBB      VDDH    VPP     VSS     h3_0    OAI22D2BM156H3P48CPDELVT_1_P_ULVTLL_L2H
x_U2_p6_3           np6_5    np4_3    VBB     VDD     VDDH    VPP     VSS     p6_3    NR2D1BM156H3P48CPDELVT_1_P_ULVTLL_L2H_V02
x_U2_h7_4           np6_5    nh5_4    nh7_6    nh7_6    VBB     VDD     VDDH    VPP     VSS     h7_4    OAI22D1BM156H3P48CPDELVT_P_ULVTLL_L2H_V02
x_U2_p10_7          np10_9    np8_7    VBB     VDD     VDDH    VPP     VSS     p10_7    NR2D1BM156H3P48CPDELVT_1_P_ULVTLL_L2H_V02
x_U2_h11_8          np10_9    nh9_8    nh11_10    nh11_10    VBB     VDD     VDDH    VPP     VSS     h11_8    OAI22D1BM156H3P48CPDELVT_P_ULVTLL_L2H_V02
x_U2_p14_11         np14_13    np12_11    VBB     VDD     VDDH    VPP     VSS     p14_11    NR2D1BM156H3P48CPDELVT_1_P_ULVTLL_L2H_V02
x_U2_h15_12         np14_13    nh13_12    nh15_14    nh15_14    VBB     VDD     VDDH    VPP     VSS     h15_12    OAI22D1BM156H3P48CPDELVT_P_ULVTLL_L2H_V02
x_U2_p18_15         np18_17    np16_15    VBB     VDD     VPP     VSS     p18_15    NR2D1BM156H3P48CPDELVT_1
x_U2_h19_16         np18_17    nh17_16    nh19_18    VBB     VDD     VPP     VSS     h19_16    OAI21D1BM156H3P48CPDELVT
x_U2_p22_19         np22_21    np20_19    VBB     VDD     VPP     VSS     p22_19    NR2D1BM156H3P48CPDELVT_1
x_U2_h23_20         np22_21    nh21_20    nh23_22    VBB     VDD     VPP     VSS     h23_20    OAI21D1BM156H3P48CPDELVT
x_U2_p26_23         np26_25    np24_23    VBB     VDD     VPP     VSS     p26_23    NR2D1BM156H3P48CPDELVT_1
x_U2_p27            np27    VBB     VDD     VPP     VSS     p27     INVD1BM156H3P48CPDELVT_1
x_U2_h27_24         np26_25    nh25_24    nh27_26    VBB     VDD     VPP     VSS     h27_24    OAI21D1BM156H3P48CPDELVT
x_U2_np29_28        nq29    np28    VBB     VDD     VPP     VSS     np29_28    OR2D1BM156H3P48CPDELVT_1
x_U3_nh7_0          p6_3    h3_0    h7_4    VBB     VDD     VDDH    VPP     VSS     nh7_0    AOI21D2BM156H3P48CPDELVT_H2H_V03
x_U3_np14_7         p14_11    p10_7    VBB     VDD     VDDH    VPP     VSS     np14_7    ND2D1BM156H3P48CPDELVT_1_H2H_V03
x_U3_nh15_8         p14_11    h11_8    h15_12    VBB     VDD     VDDH    VPP     VSS     nh15_8    AOI21D1BM156H3P48CPDELVT_H2H_V03
x_U3_np22_15        p22_19    p18_15    VBB     VDD     VPP     VSS     np22_15    ND2D1BM156H3P48CPDELVT_1
x_U3_nh23_16        p22_19    h19_16    h23_20    VBB     VDD     VPP     VSS     nh23_16    AOI21D1BM156H3P48CPDELVT
x_U3_np27_23        q27     p26_23    VBB     VDD     VPP     VSS     np27_23    ND2D1BM156H3P48CPDELVT_1
x_U3_nh28_24        a28     b28     p27     h27_24    VBB     VDD     VPP     VSS     nh28_24    AOI22D1BM156H3P48CPDELVT
x_U4_h15_0          np14_7    nh7_0    nh15_8    VBB     VDD     VDDH    VPP     VSS     h15_0    OAI21D2BM156H3P48CPDELVT_H2H_V02
x_U4_p22_15         np22_15    VBB     VDD     VPP     VSS     p22_15    INVD1BM156H3P48CPDELVT_1
x_U4_h23_16         nh23_16    VBB     VDD     VPP     VSS     h23_16    INVD1BM156H3P48CPDELVT_1
x_U4_np29_23        np29_28    np27_23    VBB     VDD     VPP     VSS     np29_23    OR2D1BM156H3P48CPDELVT_1
x_U4_ng29_24        np29_28    nh28_24    ng29    VBB     VDD     VPP     VSS     ng29_24    OA21D1BM156H3P48CPDELVT
x_U1_ng0_s0         a0      b0      ng0     VBB     VDD     VPP     VSS     s0      XNR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_np1_q1         a1      b1      np1     VBB     VDD     VPP     VSS     q1      XOR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_ng2_nq2        a2      b2      ng2     VBB     VDD     VPP     VSS     nq2     XNR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_np3_q3         a3      b3      np3     VBB     VDD     VPP     VSS     q3      XOR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_ng4_nq4        a4      b4      ng4     VBB     VDD     VPP     VSS     nq4     XNR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_np5_q5         a5      b5      np5     VBB     VDD     VPP     VSS     q5      XOR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_ng6_nq6        a6      b6      ng6     VBB     VDD     VPP     VSS     nq6     XNR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_np7_q7         a7      b7      np7     VBB     VDD     VPP     VSS     q7      XOR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_ng8_nq8        a8      b8      ng8     VBB     VDD     VPP     VSS     nq8     XNR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_np9_q9         a9      b9      np9     VBB     VDD     VPP     VSS     q9      XOR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_ng10_nq10      a10     b10     ng10    VBB     VDD     VPP     VSS     nq10    XNR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_np11_q11       a11     b11     np11    VBB     VDD     VPP     VSS     q11     XOR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_ng12_nq12      a12     b12     ng12    VBB     VDD     VPP     VSS     nq12    XNR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_np13_q13       a13     b13     np13    VBB     VDD     VPP     VSS     q13     XOR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_ng14_nq14      a14     b14     ng14    VBB     VDD     VPP     VSS     nq14    XNR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_np15_q15       a15     b15     np15    VBB     VDD     VPP     VSS     q15     XOR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_ng16_nq16      a16     b16     ng16    VBB     VDD     VPP     VSS     nq16    XNR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_np17_q17       a17     b17     np17    VBB     VDD     VPP     VSS     q17     XOR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_ng18_nq18      a18     b18     ng18    VBB     VDD     VPP     VSS     nq18    XNR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_np19_q19       a19     b19     np19    VBB     VDD     VPP     VSS     q19     XOR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_ng20_nq20      a20     b20     ng20    VBB     VDD     VPP     VSS     nq20    XNR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_np21_q21       a21     b21     np21    VBB     VDD     VPP     VSS     q21     XOR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_ng22_nq22      a22     b22     ng22    VBB     VDD     VPP     VSS     nq22    XNR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_np23_q23       a23     b23     np23    VBB     VDD     VPP     VSS     q23     XOR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_ng24_nq24      a24     b24     ng24    VBB     VDD     VPP     VSS     nq24    XNR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_np25_q25       a25     b25     np25    VBB     VDD     VPP     VSS     q25     XOR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_ng26_nq26      a26     b26     ng26    VBB     VDD     VPP     VSS     nq26    XNR2D1_DUAL_OUT_BM156H3P48CPDELVT
x_U1_nq30           a30     b30     VBB     VDD     VPP     VSS     nq30    XNR2D1BM156H3P48CPDELVT
x_U2_ng1_0          np1     nh1_0    VBB     VDD     VPP     VSS     ng1_0    OR2D1BM156H3P48CPDELVT_1
x_U2_g10_8          np10_9    nh9_8    ng10    VBB     VDD     VPP     VSS     g10_8    OAI21D1BM156H3P48CPDELVT
x_U2_g14_12         np14_13    nh13_12    ng14    VBB     VDD     VPP     VSS     g14_12    OAI21D1BM156H3P48CPDELVT
x_U2_p17_15         np17    np16_15    VBB     VDD     VPP     VSS     p17_15    NR2D1BM156H3P48CPDELVT_1
x_U2_g17_16         np17    nh17_16    VBB     VDD     VPP     VSS     g17_16    NR2D1BM156H3P48CPDELVT_1
x_U2_ng22_20        np22_21    nh21_20    ng22    VBB     VDD     VPP     VSS     ng22_20    OA21D1BM156H3P48CPDELVT
x_U2_ng26_24        np26_25    nh25_24    ng26    VBB     VDD     VPP     VSS     ng26_24    OA21D1BM156H3P48CPDELVT
x_U3_g2_0           nq2     ng1_0    ng2     VBB     VDD     VPP     VSS     g2_0    OAI21D1BM156H3P48CPDELVT
x_U3_ng3_0          np3     h3_0    VBB     VDD     VPP     VSS     ng3_0    IND2D1BM156H3P48CPDELVT_1
x_U3_np22_19        p22_19    VBB     VDD     VPP     VSS     np22_19    INVD1BM156H3P48CPDELVT_1
x_U3_np26_23        p26_23    VBB     VDD     VPP     VSS     np26_23    INVD1BM156H3P48CPDELVT_1
x_U3_ng27_24        p27     h27_24    VBB     VDD     VPP     VSS     ng27_24    ND2D1BM156H3P48CPDELVT_1
x_U4_g4_0           nq4     ng3_0    ng4     VBB     VDD     VPP     VSS     g4_0    OAI21D1BM156H3P48CPDELVT
x_U4_ng5_0          nq4     ng3_0    nh5_4    np5     VBB     VDD     VPP     VSS     ng5_0    OAO211D1BM156H3P48CPDELVT
x_U4_ng7_0          np7     nh7_0    VBB     VDD     VPP     VSS     ng7_0    OR2D1BM156H3P48CPDELVT_1
x_U4_nh11_0         p10_7    nh7_0    h11_8    VBB     VDD     VPP     VSS     nh11_0    IAOI21D1BM156H3P48CPDELVT
x_U5_g6_0           nq6     ng5_0    ng6     VBB     VDD     VPP     VSS     g6_0    OAI21D1BM156H3P48CPDELVT
x_U5_g8_0           nq8     ng7_0    ng8     VBB     VDD     VPP     VSS     g8_0    OAI21D1BM156H3P48CPDELVT
x_U5_g9_0           np8_7    ng7_0    nh9_8    np9     VBB     VDD     VPP     VSS     g9_0    OAOI211D1BM156H3P48CPDELVT
x_U5_ng10_0         p10_7    ng7_0    g10_8    VBB     VDD     VPP     VSS     ng10_0    IAOI21D1BM156H3P48CPDELVT
x_U5_g11_0          np11    nh11_0    VBB     VDD     VPP     VSS     g11_0    NR2D1BM156H3P48CPDELVT_1
x_U5_g12_0          np12_11    nh11_0    ng12    VBB     VDD     VPP     VSS     g12_0    OAI21D1BM156H3P48CPDELVT
x_U5_g13_0          np12_11    nh11_0    nh13_12    np13    VBB     VDD     VPP     VSS     g13_0    OAOI211D1BM156H3P48CPDELVT
x_U5_ng14_0         p14_11    nh11_0    g14_12    VBB     VDD     VPP     VSS     ng14_0    IAOI21D1BM156H3P48CPDELVT
x_U5_ng15_0         np15    h15_0    VBB     VDD     VPP     VSS     ng15_0    IND2D1BM156H3P48CPDELVT_1
x_U5_ng17_0         p17_15    h15_0    g17_16    VBB     VDD     VPP     VSS     ng17_0    AOI21D1BM156H3P48CPDELVT
x_U5_nh19_0         p18_15    h15_0    h19_16    VBB     VDD     VPP     VSS     nh19_0    AOI21D2BM156H3P48CPDELVT
x_U5_nh23_0         p22_15    h15_0    h23_16    VBB     VDD     VPP     VSS     nh23_0    AOI21D2BM156H3P48CPDELVT
x_U5_nh23_0_copy    p22_15    h15_0    h23_16    VBB     VDD     VPP     VSS     nh23_0    AOI21D2BM156H3P48CPDELVT
x_U6_g16_0          nq16    ng15_0    ng16    VBB     VDD     VPP     VSS     g16_0    OAI21D1BM156H3P48CPDELVT
x_U6_g18_0          nq18    ng17_0    ng18    VBB     VDD     VPP     VSS     g18_0    OAI21D1BM156H3P48CPDELVT
x_U6_g19_0          np19    nh19_0    VBB     VDD     VPP     VSS     g19_0    NR2D1BM156H3P48CPDELVT_1
x_U6_g20_0          np20_19    nh19_0    ng20    VBB     VDD     VPP     VSS     g20_0    OAI21D1BM156H3P48CPDELVT
x_U6_g21_0          np20_19    nh19_0    nh21_20    np21    VBB     VDD     VPP     VSS     g21_0    OAOI211D1BM156H3P48CPDELVT
x_U6_g22_0          np22_19    nh19_0    ng22_20    VBB     VDD     VPP     VSS     g22_0    OAI21D1BM156H3P48CPDELVT
x_U6_g23_0          np23    nh23_0    VBB     VDD     VPP     VSS     g23_0    NR2D1BM156H3P48CPDELVT_1
x_U6_g24_0          np24_23    nh23_0    ng24    VBB     VDD     VPP     VSS     g24_0    OAI21D1BM156H3P48CPDELVT
x_U6_g25_0          np24_23    nh23_0    nh25_24    np25    VBB     VDD     VPP     VSS     g25_0    OAOI211D1BM156H3P48CPDELVT
x_U6_g26_0          np26_23    nh23_0    ng26_24    VBB     VDD     VPP     VSS     g26_0    OAI21D1BM156H3P48CPDELVT
x_U6_g27_0          np27_23    nh23_0    ng27_24    VBB     VDD     VPP     VSS     g27_0    OAI21D1BM156H3P48CPDELVT
x_U6_g28_0          np27_23    nh23_0    nh28_24    np28    VBB     VDD     VPP     VSS     g28_0    OAOI211D1BM156H3P48CPDELVT
x_U6_g29_0          np29_23    nh23_0    ng29_24    VBB     VDD     VPP     VSS     g29_0    OAI21D1BM156H3P48CPDELVT
x_U2_s1             ng0     q1      VBB     VDD     VPP     VSS     s1      XOR2D1BM156H3P48CPDELVT
x_U3_s2             ng1_0    nq2     VBB     VDD     VPP     VSS     s2      XNR2D1BM156H3P48CPDELVT
x_U4_s3             g2_0    q3      VBB     VDD     VPP     VSS     s3      XNR2D1BM156H3P48CPDELVT
x_U4_s4             ng3_0    nq4     VBB     VDD     VPP     VSS     s4      XNR2D1BM156H3P48CPDELVT
x_U5_s5             g4_0    q5      VBB     VDD     VPP     VSS     s5      XNR2D1BM156H3P48CPDELVT
x_U5_s6             ng5_0    nq6     VBB     VDD     VPP     VSS     s6      XNR2D1BM156H3P48CPDELVT
x_U6_s7             g6_0    q7      VBB     VDD     VPP     VSS     s7      XNR2D1BM156H3P48CPDELVT
x_U5_s8             ng7_0    nq8     VBB     VDD     VPP     VSS     s8      XNR2D1BM156H3P48CPDELVT
x_U6_s9             g8_0    q9      VBB     VDD     VPP     VSS     s9      XNR2D1BM156H3P48CPDELVT
x_U6_s10            g9_0    nq10    VBB     VDD     VPP     VSS     s10     XOR2D1BM156H3P48CPDELVT
x_U6_s11            ng10_0    q11     VBB     VDD     VPP     VSS     s11     XOR2D1BM156H3P48CPDELVT
x_U6_s12            g11_0    nq12    VBB     VDD     VPP     VSS     s12     XOR2D1BM156H3P48CPDELVT
x_U6_s13            g12_0    q13     VBB     VDD     VPP     VSS     s13     XNR2D1BM156H3P48CPDELVT
x_U6_s14            g13_0    nq14    VBB     VDD     VPP     VSS     s14     XOR2D1BM156H3P48CPDELVT
x_U6_s15            ng14_0    q15     VBB     VDD     VPP     VSS     s15     XOR2D1BM156H3P48CPDELVT
x_U6_s16            ng15_0    nq16    VBB     VDD     VPP     VSS     s16     XNR2D1BM156H3P48CPDELVT
x_U7_s17            g16_0    q17     VBB     VDD     VPP     VSS     s17     XNR2D1BM156H3P48CPDELVT
x_U6_s18            ng17_0    nq18    VBB     VDD     VPP     VSS     s18     XNR2D1BM156H3P48CPDELVT
x_U7_s19            g18_0    q19     VBB     VDD     VPP     VSS     s19     XNR2D1BM156H3P48CPDELVT
x_U7_s20            g19_0    nq20    VBB     VDD     VPP     VSS     s20     XOR2D1BM156H3P48CPDELVT
x_U7_s21            g20_0    q21     VBB     VDD     VPP     VSS     s21     XNR2D1BM156H3P48CPDELVT
x_U7_s22            g21_0    nq22    VBB     VDD     VPP     VSS     s22     XOR2D1BM156H3P48CPDELVT
x_U7_s23            g22_0    q23     VBB     VDD     VPP     VSS     s23     XNR2D1BM156H3P48CPDELVT
x_U7_s24            g23_0    nq24    VBB     VDD     VPP     VSS     s24     XOR2D1BM156H3P48CPDELVT
x_U7_s25            g24_0    q25     VBB     VDD     VPP     VSS     s25     XNR2D1BM156H3P48CPDELVT
x_U7_s26            g25_0    nq26    VBB     VDD     VPP     VSS     s26     XOR2D1BM156H3P48CPDELVT
x_U7_s27            g26_0    q27     VBB     VDD     VPP     VSS     s27     XNR2D1BM156H3P48CPDELVT
x_U7_s28            g27_0    q28     VBB     VDD     VPP     VSS     s28     XNR2D1BM156H3P48CPDELVT
x_U7_s29            g28_0    nq29    VBB     VDD     VPP     VSS     s29     XOR2D1BM156H3P48CPDELVT
x_U7_s30            g29_0    nq30    VBB     VDD     VPP     VSS     s30     XOR2D1BM156H3P48CPDELVT
.ENDS
