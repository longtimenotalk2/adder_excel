.inc '/ic/projects/BM1340/public/5_custom/spf/stdcell/Cbest/INVMZD1BWP200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/stdcell/Cbest/ND2MZD1BWP200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/stdcell/Cbest/NR2MZD1BWP200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/stdcell/Cbest/OR2MZD1BWP200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/stdcell/Cbest/IND2NOMSAMZD1BWP200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/XOR2SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/XNR2SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/AOI21SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/AOI21SAMZD2BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/OAI21SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/OAI21SAMZD2BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/IAOI21SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/AOI22SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/OAI22SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/OAOI211SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/OAO211MZD1BM200H6P51CNODELVT.Cbest60.spf'

.SUBCKT UFADDER_PP_31_B32 A0 A1 A2 A3 A4 A5 A6 A7 A8 A9 A10 A11 A12 A13 A14 A15 A16 A17 A18 A19 A20 A21 A22 A23 A24 A25 A26 A27 A28 A29 A30 B0 B1 B2 B3 B4 B5 B6 B7 B8 B9 B10 B11 B12 B13 B14 B15 B16 B17 B18 B19 B20 B21 B22 B23 B24 B25 B26 B27 B28 B29 B30 S0 S1 S2 S3 S4 S5 S6 S7 S8 S9 S10 S11 S12 S13 S14 S15 S16 S17 S18 S19 S20 S21 S22 S23 S24 S25 S26 S27 S28 S29 S30 VBB VDD VPP VSS 
x_U1_nh1_0          a1      b1      a0      b0      VBB     VDD     VPP     VSS     nh1_0    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np2_1          a2      b2      a1      b1      VBB     VDD     VPP     VSS     np2_1    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_nh3_2          a3      b3      a2      b2      VBB     VDD     VPP     VSS     nh3_2    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np4_3          a4      b4      a3      b3      VBB     VDD     VPP     VSS     np4_3    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_nh5_4          a5      b5      a4      b4      VBB     VDD     VPP     VSS     nh5_4    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np7_6          a7      b7      a6      b6      VBB     VDD     VPP     VSS     np7_6    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_nh8_7          a8      b8      a7      b7      VBB     VDD     VPP     VSS     nh8_7    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np9_8          a9      b9      a8      b8      VBB     VDD     VPP     VSS     np9_8    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_nh10_9         a10     b10     a9      b9      VBB     VDD     VPP     VSS     nh10_9    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np11_10        a11     b11     a10     b10     VBB     VDD     VPP     VSS     np11_10    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_nh12_11        a12     b12     a11     b11     VBB     VDD     VPP     VSS     nh12_11    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np14_13        a14     b14     a13     b13     VBB     VDD     VPP     VSS     np14_13    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_nh15_14        a15     b15     a14     b14     VBB     VDD     VPP     VSS     nh15_14    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np16_15        a16     b16     a15     b15     VBB     VDD     VPP     VSS     np16_15    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_nh17_16        a17     b17     a16     b16     VBB     VDD     VPP     VSS     nh17_16    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np18_17        a18     b18     a17     b17     VBB     VDD     VPP     VSS     np18_17    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_nh19_18        a19     b19     a18     b18     VBB     VDD     VPP     VSS     nh19_18    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np20_19        a20     b20     a19     b19     VBB     VDD     VPP     VSS     np20_19    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_ng21nq21       a21     b21     ng21    VBB     VDD     VPP     VSS     nq21    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng22nq22       a22     b22     ng22    VBB     VDD     VPP     VSS     nq22    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng23           a23     b23     VBB     VDD     VPP     VSS     ng23    ND2MZD1BWP200H6P51CNODELVT
x_U1_ng24nq24       a24     b24     ng24    VBB     VDD     VPP     VSS     nq24    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np5            a5      b5      VBB     VDD     VPP     VSS     np5     NR2MZD1BWP200H6P51CNODELVT
x_U1_ng6            a6      b6      VBB     VDD     VPP     VSS     ng6     ND2MZD1BWP200H6P51CNODELVT
x_U1_np12           a12     b12     VBB     VDD     VPP     VSS     np12    NR2MZD1BWP200H6P51CNODELVT
x_U1_ng13           a13     b13     VBB     VDD     VPP     VSS     ng13    ND2MZD1BWP200H6P51CNODELVT
x_U1_ng20nq20       a20     b20     ng20    VBB     VDD     VPP     VSS     nq20    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np23q23        a23     b23     np23    VBB     VDD     VPP     VSS     q23     XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U2_h3_0           np2_1    nh1_0    nh3_2    VBB     VDD     VPP     VSS     h3_0    OAI21SAMZD2BM200H6P51CNODELVT
x_U2_p5_3           np5     np4_3    VBB     VDD     VPP     VSS     p5_3    NR2MZD1BWP200H6P51CNODELVT
x_U2_h6_4           np5     nh5_4    ng6     VBB     VDD     VPP     VSS     h6_4    OAI21SAMZD1BM200H6P51CNODELVT
x_U2_p9_6           np9_8    np7_6    VBB     VDD     VPP     VSS     p9_6    NR2MZD1BWP200H6P51CNODELVT
x_U2_h10_7          np9_8    nh8_7    nh10_9    VBB     VDD     VPP     VSS     h10_7    OAI21SAMZD1BM200H6P51CNODELVT
x_U2_p12_10         np12    np11_10    VBB     VDD     VPP     VSS     p12_10    NR2MZD1BWP200H6P51CNODELVT
x_U2_h13_11         np12    nh12_11    ng13    VBB     VDD     VPP     VSS     h13_11    OAI21SAMZD1BM200H6P51CNODELVT
x_U2_p16_13         np16_15    np14_13    VBB     VDD     VPP     VSS     p16_13    NR2MZD1BWP200H6P51CNODELVT
x_U2_h17_14         np16_15    nh15_14    nh17_16    VBB     VDD     VPP     VSS     h17_14    OAI21SAMZD1BM200H6P51CNODELVT
x_U2_p20_17         np20_19    np18_17    VBB     VDD     VPP     VSS     p20_17    NR2MZD1BWP200H6P51CNODELVT
x_U2_g20_18         np20_19    nh19_18    ng20    VBB     VDD     VPP     VSS     g20_18    OAI21SAMZD1BM200H6P51CNODELVT
x_U2_q22_21         nq22    nq21    VBB     VDD     VPP     VSS     q22_21    NR2MZD1BWP200H6P51CNODELVT
x_U2_g22_21         nq22    ng21    ng22    VBB     VDD     VPP     VSS     g22_21    OAI21SAMZD1BM200H6P51CNODELVT
x_U2_p24_23         nq24    np23    VBB     VDD     VPP     VSS     p24_23    NR2MZD1BWP200H6P51CNODELVT
x_U2_g24_23         nq24    ng23    ng24    VBB     VDD     VPP     VSS     g24_23    OAI21SAMZD1BM200H6P51CNODELVT
x_U3_nh6_0          p5_3    h3_0    h6_4    VBB     VDD     VPP     VSS     nh6_0    AOI21SAMZD2BM200H6P51CNODELVT
x_U3_np12_6         p12_10    p9_6    VBB     VDD     VPP     VSS     np12_6    ND2MZD1BWP200H6P51CNODELVT
x_U3_nh13_7         p12_10    h10_7    h13_11    VBB     VDD     VPP     VSS     nh13_7    AOI21SAMZD1BM200H6P51CNODELVT
x_U3_np20_13        p20_17    p16_13    VBB     VDD     VPP     VSS     np20_13    ND2MZD1BWP200H6P51CNODELVT
x_U3_ng20_14        p20_17    h17_14    g20_18    VBB     VDD     VPP     VSS     ng20_14    AOI21SAMZD1BM200H6P51CNODELVT
x_U3_nq24_21        p24_23    q22_21    VBB     VDD     VPP     VSS     nq24_21    ND2MZD1BWP200H6P51CNODELVT
x_U3_ng24_21        p24_23    g22_21    g24_23    VBB     VDD     VPP     VSS     ng24_21    AOI21SAMZD1BM200H6P51CNODELVT
x_U4_h13_0          np12_6    nh6_0    nh13_7    VBB     VDD     VPP     VSS     h13_0    OAI21SAMZD2BM200H6P51CNODELVT
x_U4_p24_13         nq24_21    np20_13    VBB     VDD     VPP     VSS     p24_13    NR2MZD1BWP200H6P51CNODELVT
x_U4_g24_14         nq24_21    ng20_14    ng24_21    VBB     VDD     VPP     VSS     g24_14    OAI21SAMZD1BM200H6P51CNODELVT
x_U1_ng0nq0         a0      b0      ng0     VBB     VDD     VPP     VSS     nq0     XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np1q1          a1      b1      np1     VBB     VDD     VPP     VSS     q1      XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng2nq2         a2      b2      ng2     VBB     VDD     VPP     VSS     nq2     XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np3q3          a3      b3      np3     VBB     VDD     VPP     VSS     q3      XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng4nq4         a4      b4      ng4     VBB     VDD     VPP     VSS     nq4     XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_q5             a5      b5      VBB     VDD     VPP     VSS     q5      XOR2SAMZD1BM200H6P51CNODELVT
x_U1_np6q6          a6      b6      np6     VBB     VDD     VPP     VSS     q6      XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng7nq7         a7      b7      ng7     VBB     VDD     VPP     VSS     nq7     XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np8q8          a8      b8      np8     VBB     VDD     VPP     VSS     q8      XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng9nq9         a9      b9      ng9     VBB     VDD     VPP     VSS     nq9     XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np10q10        a10     b10     np10    VBB     VDD     VPP     VSS     q10     XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng11nq11       a11     b11     ng11    VBB     VDD     VPP     VSS     nq11    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_q12            a12     b12     VBB     VDD     VPP     VSS     q12     XOR2SAMZD1BM200H6P51CNODELVT
x_U1_np13q13        a13     b13     np13    VBB     VDD     VPP     VSS     q13     XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng14nq14       a14     b14     ng14    VBB     VDD     VPP     VSS     nq14    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np15q15        a15     b15     np15    VBB     VDD     VPP     VSS     q15     XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng16nq16       a16     b16     ng16    VBB     VDD     VPP     VSS     nq16    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np17q17        a17     b17     np17    VBB     VDD     VPP     VSS     q17     XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng18nq18       a18     b18     ng18    VBB     VDD     VPP     VSS     nq18    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np19q19        a19     b19     np19    VBB     VDD     VPP     VSS     q19     XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng25nq25       a25     b25     ng25    VBB     VDD     VPP     VSS     nq25    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng26nq26       a26     b26     ng26    VBB     VDD     VPP     VSS     nq26    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_q27            a27     b27     VBB     VDD     VPP     VSS     q27     XOR2SAMZD1BM200H6P51CNODELVT
x_U1_ng28nq28       a28     b28     ng28    VBB     VDD     VPP     VSS     nq28    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_q29            a29     b29     VBB     VDD     VPP     VSS     q29     XOR2SAMZD1BM200H6P51CNODELVT
x_U1_nq30           a30     b30     VBB     VDD     VPP     VSS     nq30    XNR2SAMZD1BM200H6P51CNODELVT
x_U2_ng1_0          np1     nh1_0    VBB     VDD     VPP     VSS     ng1_0    OR2MZD1BWP200H6P51CNODELVT
x_U2_g9_7           np9_8    nh8_7    ng9     VBB     VDD     VPP     VSS     g9_7    OAI21SAMZD1BM200H6P51CNODELVT
x_U2_g16_14         np16_15    nh15_14    ng16    VBB     VDD     VPP     VSS     g16_14    OAI21SAMZD1BM200H6P51CNODELVT
x_U2_nq23_21        q23     q22_21    VBB     VDD     VPP     VSS     nq23_21    ND2MZD1BWP200H6P51CNODELVT
x_U2_ng23_21        a23     b23     q23     g22_21    VBB     VDD     VPP     VSS     ng23_21    AOI22SAMZD1BM200H6P51CNODELVT
x_U2_q26_25         nq26    nq25    VBB     VDD     VPP     VSS     q26_25    NR2MZD1BWP200H6P51CNODELVT
x_U2_g26_25         nq26    ng25    ng26    VBB     VDD     VPP     VSS     g26_25    OAI21SAMZD1BM200H6P51CNODELVT
x_U3_g2_0           nq2     ng1_0    ng2     VBB     VDD     VPP     VSS     g2_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U3_ng3_0          np3     h3_0    VBB     VDD     VPP     VSS     ng3_0    IND2NOMSAMZD1BWP200H6P51CNODELVT
x_U3_nq22_21        q22_21    VBB     VDD     VPP     VSS     nq22_21    INVMZD1BWP200H6P51CNODELVT
x_U3_ng22_21        g22_21    VBB     VDD     VPP     VSS     ng22_21    INVMZD1BWP200H6P51CNODELVT
x_U3_nq27_25        q27     q26_25    VBB     VDD     VPP     VSS     nq27_25    ND2MZD1BWP200H6P51CNODELVT
x_U3_ng27_25        a27     b27     q27     g26_25    VBB     VDD     VPP     VSS     ng27_25    AOI22SAMZD1BM200H6P51CNODELVT
x_U4_g4_0           nq4     ng3_0    ng4     VBB     VDD     VPP     VSS     g4_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U4_ng5_0          ng3_0    nq4     nh5_4    np5     VBB     VDD     VPP     VSS     ng5_0    OAO211MZD1BM200H6P51CNODELVT
x_U4_ng6_0          np6     nh6_0    VBB     VDD     VPP     VSS     ng6_0    OR2MZD1BWP200H6P51CNODELVT
x_U4_nh10_0         p9_6    nh6_0    h10_7    VBB     VDD     VPP     VSS     nh10_0    IAOI21SAMZD1BM200H6P51CNODELVT
x_U4_p20_13         np20_13    VBB     VDD     VPP     VSS     p20_13    INVMZD1BWP200H6P51CNODELVT
x_U4_g20_14         ng20_14    VBB     VDD     VPP     VSS     g20_14    INVMZD1BWP200H6P51CNODELVT
x_U4_q28_25         nq28    nq27_25    VBB     VDD     VPP     VSS     q28_25    NR2MZD1BWP200H6P51CNODELVT
x_U4_g28_25         nq28    ng27_25    ng28    VBB     VDD     VPP     VSS     g28_25    OAI21SAMZD1BM200H6P51CNODELVT
x_U5_g7_0           nq7     ng6_0    ng7     VBB     VDD     VPP     VSS     g7_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U5_g8_0           ng6_0    np7_6    nh8_7    np8     VBB     VDD     VPP     VSS     g8_0    OAOI211SAMZD1BM200H6P51CNODELVT
x_U5_ng9_0          p9_6    ng6_0    g9_7    VBB     VDD     VPP     VSS     ng9_0    IAOI21SAMZD1BM200H6P51CNODELVT
x_U5_g10_0          np10    nh10_0    VBB     VDD     VPP     VSS     g10_0    NR2MZD1BWP200H6P51CNODELVT
x_U5_g11_0          np11_10    nh10_0    ng11    VBB     VDD     VPP     VSS     g11_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U5_g12_0          nh10_0    np11_10    nh12_11    np12    VBB     VDD     VPP     VSS     g12_0    OAOI211SAMZD1BM200H6P51CNODELVT
x_U5_nh13_0         h13_0    VBB     VDD     VPP     VSS     nh13_0    INVMZD1BWP200H6P51CNODELVT
x_U5_nh17_0         p16_13    h13_0    h17_14    VBB     VDD     VPP     VSS     nh17_0    AOI21SAMZD1BM200H6P51CNODELVT
x_U5_ng20_0         p20_13    h13_0    g20_14    VBB     VDD     VPP     VSS     ng20_0    AOI21SAMZD1BM200H6P51CNODELVT
x_U5_ng24_0         p24_13    h13_0    g24_14    VBB     VDD     VPP     VSS     ng24_0    AOI21SAMZD2BM200H6P51CNODELVT
x_U5_nq29_25        q29     q28_25    VBB     VDD     VPP     VSS     nq29_25    ND2MZD1BWP200H6P51CNODELVT
x_U5_ng29_25        a29     b29     q29     g28_25    VBB     VDD     VPP     VSS     ng29_25    AOI22SAMZD1BM200H6P51CNODELVT
x_U6_g13_0          np13    nh13_0    VBB     VDD     VPP     VSS     g13_0    NR2MZD1BWP200H6P51CNODELVT
x_U6_g14_0          np14_13    nh13_0    ng14    VBB     VDD     VPP     VSS     g14_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g15_0          nh13_0    np14_13    nh15_14    np15    VBB     VDD     VPP     VSS     g15_0    OAOI211SAMZD1BM200H6P51CNODELVT
x_U6_ng16_0         p16_13    nh13_0    g16_14    VBB     VDD     VPP     VSS     ng16_0    IAOI21SAMZD1BM200H6P51CNODELVT
x_U6_g17_0          np17    nh17_0    VBB     VDD     VPP     VSS     g17_0    NR2MZD1BWP200H6P51CNODELVT
x_U6_g18_0          np18_17    nh17_0    ng18    VBB     VDD     VPP     VSS     g18_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g19_0          nh17_0    np18_17    nh19_18    np19    VBB     VDD     VPP     VSS     g19_0    OAOI211SAMZD1BM200H6P51CNODELVT
x_U6_g21_0          nq21    ng20_0    ng21    VBB     VDD     VPP     VSS     g21_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g22_0          nq22_21    ng20_0    ng22_21    VBB     VDD     VPP     VSS     g22_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g23_0          nq23_21    ng20_0    ng23_21    VBB     VDD     VPP     VSS     g23_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g24_0          ng24_0    VBB     VDD     VPP     VSS     g24_0    INVMZD1BWP200H6P51CNODELVT
x_U6_g25_0          nq25    ng24_0    ng25    VBB     VDD     VPP     VSS     g25_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g27_0          nq27_25    ng24_0    ng27_25    VBB     VDD     VPP     VSS     g27_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g29_0          nq29_25    ng24_0    ng29_25    VBB     VDD     VPP     VSS     g29_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U7_ng26_0         q26_25    g24_0    g26_25    VBB     VDD     VPP     VSS     ng26_0    AOI21SAMZD1BM200H6P51CNODELVT
x_U7_ng28_0         q28_25    g24_0    g28_25    VBB     VDD     VPP     VSS     ng28_0    AOI21SAMZD1BM200H6P51CNODELVT
x_U10_s0            nq0     VBB     VDD     VPP     VSS     s0      INVMZD1BWP200H6P51CNODELVT
x_U10_s1            ng0     q1      VBB     VDD     VPP     VSS     s1      XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s2            ng1_0    nq2     VBB     VDD     VPP     VSS     s2      XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s3            g2_0    q3      VBB     VDD     VPP     VSS     s3      XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s4            ng3_0    nq4     VBB     VDD     VPP     VSS     s4      XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s5            g4_0    q5      VBB     VDD     VPP     VSS     s5      XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s6            ng5_0    q6      VBB     VDD     VPP     VSS     s6      XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s7            ng6_0    nq7     VBB     VDD     VPP     VSS     s7      XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s8            g7_0    q8      VBB     VDD     VPP     VSS     s8      XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s9            g8_0    nq9     VBB     VDD     VPP     VSS     s9      XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s10           ng9_0    q10     VBB     VDD     VPP     VSS     s10     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s11           g10_0    nq11    VBB     VDD     VPP     VSS     s11     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s12           g11_0    q12     VBB     VDD     VPP     VSS     s12     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s13           g12_0    q13     VBB     VDD     VPP     VSS     s13     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s14           g13_0    nq14    VBB     VDD     VPP     VSS     s14     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s15           g14_0    q15     VBB     VDD     VPP     VSS     s15     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s16           g15_0    nq16    VBB     VDD     VPP     VSS     s16     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s17           ng16_0    q17     VBB     VDD     VPP     VSS     s17     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s18           g17_0    nq18    VBB     VDD     VPP     VSS     s18     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s19           g18_0    q19     VBB     VDD     VPP     VSS     s19     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s20           g19_0    nq20    VBB     VDD     VPP     VSS     s20     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s21           ng20_0    nq21    VBB     VDD     VPP     VSS     s21     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s22           g21_0    nq22    VBB     VDD     VPP     VSS     s22     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s23           g22_0    q23     VBB     VDD     VPP     VSS     s23     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s24           g23_0    nq24    VBB     VDD     VPP     VSS     s24     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s25           g24_0    nq25    VBB     VDD     VPP     VSS     s25     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s26           g25_0    nq26    VBB     VDD     VPP     VSS     s26     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s27           ng26_0    q27     VBB     VDD     VPP     VSS     s27     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s28           g27_0    nq28    VBB     VDD     VPP     VSS     s28     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s29           ng28_0    q29     VBB     VDD     VPP     VSS     s29     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s30           g29_0    nq30    VBB     VDD     VPP     VSS     s30     XNR2SAMZD1BM200H6P51CNODELVT
.ENDS
