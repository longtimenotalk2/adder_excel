.inc '/ic/projects/BM1340/public/5_custom/spf/stdcell/Cbest/INVMZD1BWP200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/stdcell/Cbest/ND2MZD1BWP200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/stdcell/Cbest/NR2MZD1BWP200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/stdcell/Cbest/OR2MZD1BWP200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/stdcell/Cbest/IND2NOMSAMZD1BWP200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/XOR2SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/XNR2SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/AOI21SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/AOI21SAMZD2BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/OAI21SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/OAI21SAMZD2BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/OA21SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/IAOI21SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/AOI22SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/OAI22SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/OAOI211SAMZD1BM200H6P51CNODELVT.Cbest60.spf'
.inc '/ic/projects/BM1340/public/5_custom/spf/custom/Cbest/OAO211MZD1BM200H6P51CNODELVT.Cbest60.spf'

.SUBCKT UFADDER_PP_31_BASE_10 A0 A1 A2 A3 A4 A5 A6 A7 A8 A9 A10 A11 A12 A13 A14 A15 A16 A17 A18 A19 A20 A21 A22 A23 A24 A25 A26 A27 A28 A29 A30 B0 B1 B2 B3 B4 B5 B6 B7 B8 B9 B10 B11 B12 B13 B14 B15 B16 B17 B18 B19 B20 B21 B22 B23 B24 B25 B26 B27 B28 B29 B30 S0 S1 S2 S3 S4 S5 S6 S7 S8 S9 S10 S11 S12 S13 S14 S15 S16 S17 S18 S19 S20 S21 S22 S23 S24 S25 S26 S27 S28 S29 S30 VBB VDD VPP VSS 
x_U1_nh1_0          a1      b1      a0      b0      VBB     VDD     VPP     VSS     nh1_0    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np2_1          a2      b2      a1      b1      VBB     VDD     VPP     VSS     np2_1    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_nh3_2          a3      b3      a2      b2      VBB     VDD     VPP     VSS     nh3_2    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np4_3          a4      b4      a3      b3      VBB     VDD     VPP     VSS     np4_3    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_nh5_4          a5      b5      a4      b4      VBB     VDD     VPP     VSS     nh5_4    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np6_5          a6      b6      a5      b5      VBB     VDD     VPP     VSS     np6_5    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_nh7_6          a7      b7      a6      b6      VBB     VDD     VPP     VSS     nh7_6    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np8_7          a8      b8      a7      b7      VBB     VDD     VPP     VSS     np8_7    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_nh9_8          a9      b9      a8      b8      VBB     VDD     VPP     VSS     nh9_8    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np10_9         a10     b10     a9      b9      VBB     VDD     VPP     VSS     np10_9    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_nh11_10        a11     b11     a10     b10     VBB     VDD     VPP     VSS     nh11_10    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np12_11        a12     b12     a11     b11     VBB     VDD     VPP     VSS     np12_11    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_nh13_12        a13     b13     a12     b12     VBB     VDD     VPP     VSS     nh13_12    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np14_13        a14     b14     a13     b13     VBB     VDD     VPP     VSS     np14_13    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_nh15_14        a15     b15     a14     b14     VBB     VDD     VPP     VSS     nh15_14    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np16_15        a16     b16     a15     b15     VBB     VDD     VPP     VSS     np16_15    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_nh17_16        a17     b17     a16     b16     VBB     VDD     VPP     VSS     nh17_16    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np18_17        a18     b18     a17     b17     VBB     VDD     VPP     VSS     np18_17    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_np19           a19     b19     VBB     VDD     VPP     VSS     np19    NR2MZD1BWP200H6P51CNODELVT
x_U1_nh20_19        a20     b20     a19     b19     VBB     VDD     VPP     VSS     nh20_19    AOI22SAMZD1BM200H6P51CNODELVT
x_U1_np21_20        a21     b21     a20     b20     VBB     VDD     VPP     VSS     np21_20    OAI22SAMZD1BM200H6P51CNODELVT
x_U1_ng22nq22       a22     b22     ng22    VBB     VDD     VPP     VSS     nq22    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng23nq23       a23     b23     ng23    VBB     VDD     VPP     VSS     nq23    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np24q24        a24     b24     np24    VBB     VDD     VPP     VSS     q24     XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng18nq18       a18     b18     ng18    VBB     VDD     VPP     VSS     nq18    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng21nq21       a21     b21     ng21    VBB     VDD     VPP     VSS     nq21    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U2_h3_0           np2_1    nh1_0    nh3_2    VBB     VDD     VPP     VSS     h3_0    OAI21SAMZD2BM200H6P51CNODELVT
x_U2_p6_3           np6_5    np4_3    VBB     VDD     VPP     VSS     p6_3    NR2MZD1BWP200H6P51CNODELVT
x_U2_h7_4           np6_5    nh5_4    nh7_6    VBB     VDD     VPP     VSS     h7_4    OAI21SAMZD1BM200H6P51CNODELVT
x_U2_p10_7          np10_9    np8_7    VBB     VDD     VPP     VSS     p10_7    NR2MZD1BWP200H6P51CNODELVT
x_U2_h11_8          np10_9    nh9_8    nh11_10    VBB     VDD     VPP     VSS     h11_8    OAI21SAMZD1BM200H6P51CNODELVT
x_U2_p14_11         np14_13    np12_11    VBB     VDD     VPP     VSS     p14_11    NR2MZD1BWP200H6P51CNODELVT
x_U2_h15_12         np14_13    nh13_12    nh15_14    VBB     VDD     VPP     VSS     h15_12    OAI21SAMZD1BM200H6P51CNODELVT
x_U2_p18_15         np18_17    np16_15    VBB     VDD     VPP     VSS     p18_15    NR2MZD1BWP200H6P51CNODELVT
x_U2_g18_16         np18_17    nh17_16    ng18    VBB     VDD     VPP     VSS     g18_16    OAI21SAMZD1BM200H6P51CNODELVT
x_U2_p21_19         np21_20    np19    VBB     VDD     VPP     VSS     p21_19    NR2MZD1BWP200H6P51CNODELVT
x_U2_g21_19         np21_20    nh20_19    ng21    VBB     VDD     VPP     VSS     g21_19    OAI21SAMZD1BM200H6P51CNODELVT
x_U2_q23_22         nq23    nq22    VBB     VDD     VPP     VSS     q23_22    NR2MZD1BWP200H6P51CNODELVT
x_U2_g23_22         nq23    ng22    ng23    VBB     VDD     VPP     VSS     g23_22    OAI21SAMZD1BM200H6P51CNODELVT
x_U3_nh7_0          p6_3    h3_0    h7_4    VBB     VDD     VPP     VSS     nh7_0    AOI21SAMZD2BM200H6P51CNODELVT
x_U3_np14_7         p14_11    p10_7    VBB     VDD     VPP     VSS     np14_7    ND2MZD1BWP200H6P51CNODELVT
x_U3_nh15_8         p14_11    h11_8    h15_12    VBB     VDD     VPP     VSS     nh15_8    AOI21SAMZD1BM200H6P51CNODELVT
x_U3_np21_15        p21_19    p18_15    VBB     VDD     VPP     VSS     np21_15    ND2MZD1BWP200H6P51CNODELVT
x_U3_ng21_16        p21_19    g18_16    g21_19    VBB     VDD     VPP     VSS     ng21_16    AOI21SAMZD1BM200H6P51CNODELVT
x_U3_nq24_22        q24     q23_22    VBB     VDD     VPP     VSS     nq24_22    ND2MZD1BWP200H6P51CNODELVT
x_U3_ng24_22        a24     b24     q24     g23_22    VBB     VDD     VPP     VSS     ng24_22    AOI22SAMZD1BM200H6P51CNODELVT
x_U4_h15_0          np14_7    nh7_0    nh15_8    VBB     VDD     VPP     VSS     h15_0    OAI21SAMZD2BM200H6P51CNODELVT
x_U4_p24_15         nq24_22    np21_15    VBB     VDD     VPP     VSS     p24_15    NR2MZD1BWP200H6P51CNODELVT
x_U4_g24_16         nq24_22    ng21_16    ng24_22    VBB     VDD     VPP     VSS     g24_16    OAI21SAMZD1BM200H6P51CNODELVT
x_U1_ng0nq0         a0      b0      ng0     VBB     VDD     VPP     VSS     nq0     XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np1q1          a1      b1      np1     VBB     VDD     VPP     VSS     q1      XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng2nq2         a2      b2      ng2     VBB     VDD     VPP     VSS     nq2     XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np3q3          a3      b3      np3     VBB     VDD     VPP     VSS     q3      XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng4nq4         a4      b4      ng4     VBB     VDD     VPP     VSS     nq4     XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng5nq5         a5      b5      ng5     VBB     VDD     VPP     VSS     nq5     XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng6nq6         a6      b6      ng6     VBB     VDD     VPP     VSS     nq6     XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np7q7          a7      b7      np7     VBB     VDD     VPP     VSS     q7      XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng8nq8         a8      b8      ng8     VBB     VDD     VPP     VSS     nq8     XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np9q9          a9      b9      np9     VBB     VDD     VPP     VSS     q9      XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng10nq10       a10     b10     ng10    VBB     VDD     VPP     VSS     nq10    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np11q11        a11     b11     np11    VBB     VDD     VPP     VSS     q11     XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng12nq12       a12     b12     ng12    VBB     VDD     VPP     VSS     nq12    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np13q13        a13     b13     np13    VBB     VDD     VPP     VSS     q13     XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng14nq14       a14     b14     ng14    VBB     VDD     VPP     VSS     nq14    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np15q15        a15     b15     np15    VBB     VDD     VPP     VSS     q15     XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng16nq16       a16     b16     ng16    VBB     VDD     VPP     VSS     nq16    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np17q17        a17     b17     np17    VBB     VDD     VPP     VSS     q17     XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng19nq19       a19     b19     ng19    VBB     VDD     VPP     VSS     nq19    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_np20q20        a20     b20     np20    VBB     VDD     VPP     VSS     q20     XOR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng25nq25       a25     b25     ng25    VBB     VDD     VPP     VSS     nq25    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_ng26nq26       a26     b26     ng26    VBB     VDD     VPP     VSS     nq26    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_q27            a27     b27     VBB     VDD     VPP     VSS     q27     XOR2SAMZD1BM200H6P51CNODELVT
x_U1_ng28nq28       a28     b28     ng28    VBB     VDD     VPP     VSS     nq28    XNR2SAMZD1_DUAL_OUT_BM200H6P51CNODELVT
x_U1_q29            a29     b29     VBB     VDD     VPP     VSS     q29     XOR2SAMZD1BM200H6P51CNODELVT
x_U1_nq30           a30     b30     VBB     VDD     VPP     VSS     nq30    XNR2SAMZD1BM200H6P51CNODELVT
x_U2_ng1_0          np1     nh1_0    VBB     VDD     VPP     VSS     ng1_0    OR2MZD1BWP200H6P51CNODELVT
x_U2_p15            np15    VBB     VDD     VPP     VSS     p15     INVMZD1BWP200H6P51CNODELVT
x_U2_q26_25         nq26    nq25    VBB     VDD     VPP     VSS     q26_25    NR2MZD1BWP200H6P51CNODELVT
x_U2_g26_25         nq26    ng25    ng26    VBB     VDD     VPP     VSS     g26_25    OAI21SAMZD1BM200H6P51CNODELVT
x_U3_g2_0           nq2     ng1_0    ng2     VBB     VDD     VPP     VSS     g2_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U3_ng3_0          np3     h3_0    VBB     VDD     VPP     VSS     ng3_0    IND2NOMSAMZD1BWP200H6P51CNODELVT
x_U3_nq27_25        q27     q26_25    VBB     VDD     VPP     VSS     nq27_25    ND2MZD1BWP200H6P51CNODELVT
x_U3_ng27_25        a27     b27     q27     g26_25    VBB     VDD     VPP     VSS     ng27_25    AOI22SAMZD1BM200H6P51CNODELVT
x_U3_nq23_22        q23_22    VBB     VDD     VPP     VSS     nq23_22    INVMZD1BWP200H6P51CNODELVT
x_U3_ng23_22        g23_22    VBB     VDD     VPP     VSS     ng23_22    INVMZD1BWP200H6P51CNODELVT
x_U4_ng4_0          nq4     ng3_0    ng4     VBB     VDD     VPP     VSS     ng4_0    OA21SAMZD1BM200H6P51CNODELVT
x_U4_ng7_0          np7     nh7_0    VBB     VDD     VPP     VSS     ng7_0    OR2MZD1BWP200H6P51CNODELVT
x_U4_nh11_0         p10_7    nh7_0    h11_8    VBB     VDD     VPP     VSS     nh11_0    IAOI21SAMZD1BM200H6P51CNODELVT
x_U4_p21_15         np21_15    VBB     VDD     VPP     VSS     p21_15    INVMZD1BWP200H6P51CNODELVT
x_U4_g21_16         ng21_16    VBB     VDD     VPP     VSS     g21_16    INVMZD1BWP200H6P51CNODELVT
x_U4_q28_25         nq28    nq27_25    VBB     VDD     VPP     VSS     q28_25    NR2MZD1BWP200H6P51CNODELVT
x_U4_g28_25         nq28    ng27_25    ng28    VBB     VDD     VPP     VSS     g28_25    OAI21SAMZD1BM200H6P51CNODELVT
x_U5_ng5_0          nq5     ng4_0    ng5     VBB     VDD     VPP     VSS     ng5_0    OA21SAMZD1BM200H6P51CNODELVT
x_U5_g8_0           nq8     ng7_0    ng8     VBB     VDD     VPP     VSS     g8_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U5_ng9_0          ng7_0    np8_7    nh9_8    np9     VBB     VDD     VPP     VSS     ng9_0    OAO211MZD1BM200H6P51CNODELVT
x_U5_ng11_0         np11    nh11_0    VBB     VDD     VPP     VSS     ng11_0    OR2MZD1BWP200H6P51CNODELVT
x_U5_ng13_0         nh11_0    np12_11    nh13_12    np13    VBB     VDD     VPP     VSS     ng13_0    OAO211MZD1BM200H6P51CNODELVT
x_U5_ng15_0         p15     h15_0    VBB     VDD     VPP     VSS     ng15_0    ND2MZD1BWP200H6P51CNODELVT
x_U5_ng18_0         p18_15    h15_0    g18_16    VBB     VDD     VPP     VSS     ng18_0    AOI21SAMZD1BM200H6P51CNODELVT
x_U5_ng21_0         p21_15    h15_0    g21_16    VBB     VDD     VPP     VSS     ng21_0    AOI21SAMZD1BM200H6P51CNODELVT
x_U5_ng24_0         p24_15    h15_0    g24_16    VBB     VDD     VPP     VSS     ng24_0    AOI21SAMZD2BM200H6P51CNODELVT
x_U5_nq29_25        q29     q28_25    VBB     VDD     VPP     VSS     nq29_25    ND2MZD1BWP200H6P51CNODELVT
x_U5_ng29_25        a29     b29     q29     g28_25    VBB     VDD     VPP     VSS     ng29_25    AOI22SAMZD1BM200H6P51CNODELVT
x_U6_g6_0           nq6     ng5_0    ng6     VBB     VDD     VPP     VSS     g6_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g10_0          nq10    ng9_0    ng10    VBB     VDD     VPP     VSS     g10_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g12_0          nq12    ng11_0    ng12    VBB     VDD     VPP     VSS     g12_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g14_0          nq14    ng13_0    ng14    VBB     VDD     VPP     VSS     g14_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g16_0          nq16    ng15_0    ng16    VBB     VDD     VPP     VSS     g16_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g17_0          ng15_0    nq16    nh17_16    np17    VBB     VDD     VPP     VSS     g17_0    OAOI211SAMZD1BM200H6P51CNODELVT
x_U6_g19_0          nq19    ng18_0    ng19    VBB     VDD     VPP     VSS     g19_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g20_0          ng18_0    nq19    nh20_19    np20    VBB     VDD     VPP     VSS     g20_0    OAOI211SAMZD1BM200H6P51CNODELVT
x_U6_g22_0          nq22    ng21_0    ng22    VBB     VDD     VPP     VSS     g22_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g23_0          nq23_22    ng21_0    ng23_22    VBB     VDD     VPP     VSS     g23_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g24_0          ng24_0    VBB     VDD     VPP     VSS     g24_0    INVMZD1BWP200H6P51CNODELVT
x_U6_g25_0          nq25    ng24_0    ng25    VBB     VDD     VPP     VSS     g25_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g27_0          nq27_25    ng24_0    ng27_25    VBB     VDD     VPP     VSS     g27_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U6_g29_0          nq29_25    ng24_0    ng29_25    VBB     VDD     VPP     VSS     g29_0    OAI21SAMZD1BM200H6P51CNODELVT
x_U7_ng26_0         q26_25    g24_0    g26_25    VBB     VDD     VPP     VSS     ng26_0    AOI21SAMZD1BM200H6P51CNODELVT
x_U7_ng28_0         q28_25    g24_0    g28_25    VBB     VDD     VPP     VSS     ng28_0    AOI21SAMZD1BM200H6P51CNODELVT
x_U10_s0            nq0     VBB     VDD     VPP     VSS     s0      INVMZD1BWP200H6P51CNODELVT
x_U10_s1            ng0     q1      VBB     VDD     VPP     VSS     s1      XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s2            ng1_0    nq2     VBB     VDD     VPP     VSS     s2      XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s3            g2_0    q3      VBB     VDD     VPP     VSS     s3      XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s4            ng3_0    nq4     VBB     VDD     VPP     VSS     s4      XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s5            ng4_0    nq5     VBB     VDD     VPP     VSS     s5      XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s6            ng5_0    nq6     VBB     VDD     VPP     VSS     s6      XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s7            g6_0    q7      VBB     VDD     VPP     VSS     s7      XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s8            ng7_0    nq8     VBB     VDD     VPP     VSS     s8      XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s9            g8_0    q9      VBB     VDD     VPP     VSS     s9      XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s10           ng9_0    nq10    VBB     VDD     VPP     VSS     s10     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s11           g10_0    q11     VBB     VDD     VPP     VSS     s11     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s12           ng11_0    nq12    VBB     VDD     VPP     VSS     s12     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s13           g12_0    q13     VBB     VDD     VPP     VSS     s13     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s14           ng13_0    nq14    VBB     VDD     VPP     VSS     s14     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s15           g14_0    q15     VBB     VDD     VPP     VSS     s15     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s16           ng15_0    nq16    VBB     VDD     VPP     VSS     s16     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s17           g16_0    q17     VBB     VDD     VPP     VSS     s17     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s18           g17_0    nq18    VBB     VDD     VPP     VSS     s18     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s19           ng18_0    nq19    VBB     VDD     VPP     VSS     s19     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s20           g19_0    q20     VBB     VDD     VPP     VSS     s20     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s21           g20_0    nq21    VBB     VDD     VPP     VSS     s21     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s22           ng21_0    nq22    VBB     VDD     VPP     VSS     s22     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s23           g22_0    nq23    VBB     VDD     VPP     VSS     s23     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s24           g23_0    q24     VBB     VDD     VPP     VSS     s24     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s25           ng24_0    nq25    VBB     VDD     VPP     VSS     s25     XOR2SAMZD1BM200H6P51CNODELVT
x_U10_s26           g25_0    nq26    VBB     VDD     VPP     VSS     s26     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s27           ng26_0    q27     VBB     VDD     VPP     VSS     s27     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s28           g27_0    nq28    VBB     VDD     VPP     VSS     s28     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s29           ng28_0    q29     VBB     VDD     VPP     VSS     s29     XNR2SAMZD1BM200H6P51CNODELVT
x_U10_s30           g29_0    nq30    VBB     VDD     VPP     VSS     s30     XNR2SAMZD1BM200H6P51CNODELVT
.ENDS
